module src

struct Article {
	id		   	int
	created_at 	int
mut:
	author		string
	project 	string
	name 		string
	description string
	url			string
}
