module src

pub fn (mut app App) add_profile(profile Profile) {

	// println( app.db.exec("select full_name from profiles where full_name=$profile.full_name")[0] )

	// if full_name_len == 0 {
	// 	sql app.db {
	// 		insert profile into Profile
	// 	}
	// }
}