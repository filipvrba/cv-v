module src

struct AdminLoggedIn {
	admin_token  string
	admin_logout int
}
