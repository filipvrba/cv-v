module src

struct Profile {
	id		   int
	created_at int
mut:
	full_name string
	avatar	  string
	email     string
	phone	  string
	bio		  string
}